`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:06:11 02/28/2022 
// Design Name: 
// Module Name:    Mux4to1_LM_19101664 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Mux4to1_LM_19101664(
    input I0,
    input I1,
    input I2,
    input I3,
    input S0,
    input S1
    );


endmodule
